library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity Slave is
	
	Port (
		i_CLK		: std_logic
	);
end Slave;